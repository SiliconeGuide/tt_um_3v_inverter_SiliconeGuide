magic
tech sky130A
magscale 1 2
timestamp 1757259024
<< viali >>
rect 3822 28 4036 64
rect 5994 0 9208 40
rect 3782 -2288 4010 -2248
rect 5978 -2266 9212 -2226
<< metal1 >>
rect 3222 830 9942 1030
rect 3222 -120 3422 830
rect 3806 514 9222 830
rect 3806 64 4046 514
rect 3806 28 3822 64
rect 4036 28 4046 64
rect 3806 12 4046 28
rect 5982 40 9222 514
rect 5982 0 5994 40
rect 9208 0 9222 40
rect 5982 -10 9222 0
rect 4532 -120 5242 -118
rect 9719 -120 9801 830
rect 3222 -260 3862 -120
rect 3222 -266 3422 -260
rect 3978 -264 5242 -120
rect 5988 -188 5998 -134
rect 6052 -188 6062 -134
rect 6304 -188 6314 -134
rect 6368 -188 6378 -134
rect 6620 -188 6630 -134
rect 6684 -188 6694 -134
rect 6936 -188 6946 -134
rect 7000 -188 7010 -134
rect 7252 -188 7262 -134
rect 7316 -188 7326 -134
rect 7568 -188 7578 -134
rect 7632 -188 7642 -134
rect 7884 -188 7894 -134
rect 7948 -188 7958 -134
rect 8200 -188 8210 -134
rect 8264 -188 8274 -134
rect 8516 -188 8526 -134
rect 8580 -188 8590 -134
rect 8832 -188 8842 -134
rect 8896 -188 8906 -134
rect 9148 -188 9158 -134
rect 9212 -188 9222 -134
rect 9713 -202 9719 -120
rect 9801 -202 9807 -120
rect 2992 -382 3976 -334
rect 4532 -360 5242 -264
rect 6144 -304 6154 -250
rect 6208 -304 6218 -250
rect 6460 -304 6470 -250
rect 6524 -304 6534 -250
rect 6776 -304 6786 -250
rect 6840 -304 6850 -250
rect 7092 -304 7102 -250
rect 7156 -304 7166 -250
rect 7408 -304 7418 -250
rect 7472 -304 7482 -250
rect 7724 -304 7734 -250
rect 7788 -304 7798 -250
rect 8040 -304 8050 -250
rect 8104 -304 8114 -250
rect 8356 -304 8366 -250
rect 8420 -304 8430 -250
rect 8672 -304 8682 -250
rect 8736 -304 8746 -250
rect 8988 -304 8998 -250
rect 9052 -304 9062 -250
rect 9841 -318 9847 -236
rect 9929 -318 9935 -236
rect 2992 -1848 3192 -382
rect 4532 -408 9158 -360
rect 4532 -1828 5242 -408
rect 9847 -982 9929 -318
rect 9784 -1182 9984 -982
rect 2992 -1896 3944 -1848
rect 4532 -1876 9150 -1828
rect 3232 -1956 3432 -1950
rect 3232 -2100 3832 -1956
rect 4532 -1958 5242 -1876
rect 9847 -1900 9937 -1182
rect 3232 -2830 3432 -2100
rect 3950 -2102 5242 -1958
rect 5978 -1976 5988 -1922
rect 6042 -1976 6052 -1922
rect 6294 -1976 6304 -1922
rect 6358 -1976 6368 -1922
rect 6610 -1976 6620 -1922
rect 6674 -1976 6684 -1922
rect 6926 -1976 6936 -1922
rect 6990 -1976 7000 -1922
rect 7242 -1976 7252 -1922
rect 7306 -1976 7316 -1922
rect 7558 -1976 7568 -1922
rect 7622 -1976 7632 -1922
rect 7874 -1976 7884 -1922
rect 7938 -1976 7948 -1922
rect 8190 -1976 8200 -1922
rect 8254 -1976 8264 -1922
rect 8506 -1976 8516 -1922
rect 8570 -1976 8580 -1922
rect 8822 -1976 8832 -1922
rect 8886 -1976 8896 -1922
rect 9138 -1976 9148 -1922
rect 9202 -1976 9212 -1922
rect 9841 -1990 9847 -1900
rect 9937 -1990 9943 -1900
rect 6134 -2090 6144 -2036
rect 6198 -2090 6208 -2036
rect 6450 -2090 6460 -2036
rect 6514 -2090 6524 -2036
rect 6766 -2090 6776 -2036
rect 6830 -2090 6840 -2036
rect 7082 -2090 7092 -2036
rect 7146 -2090 7156 -2036
rect 7398 -2090 7408 -2036
rect 7462 -2090 7472 -2036
rect 7714 -2090 7724 -2036
rect 7778 -2090 7788 -2036
rect 8030 -2090 8040 -2036
rect 8094 -2090 8104 -2036
rect 8346 -2090 8356 -2036
rect 8410 -2090 8420 -2036
rect 8662 -2090 8672 -2036
rect 8726 -2090 8736 -2036
rect 8978 -2090 8988 -2036
rect 9042 -2090 9052 -2036
rect 5966 -2226 9224 -2212
rect 3764 -2248 4020 -2236
rect 3764 -2288 3782 -2248
rect 4010 -2288 4020 -2248
rect 3764 -2548 4020 -2288
rect 5966 -2266 5978 -2226
rect 9212 -2266 9224 -2226
rect 9601 -2253 9607 -2171
rect 9689 -2253 9695 -2171
rect 5966 -2548 9224 -2266
rect 3764 -2830 9224 -2548
rect 9607 -2830 9689 -2253
rect 3232 -3030 9934 -2830
<< via1 >>
rect 5998 -188 6052 -134
rect 6314 -188 6368 -134
rect 6630 -188 6684 -134
rect 6946 -188 7000 -134
rect 7262 -188 7316 -134
rect 7578 -188 7632 -134
rect 7894 -188 7948 -134
rect 8210 -188 8264 -134
rect 8526 -188 8580 -134
rect 8842 -188 8896 -134
rect 9158 -188 9212 -134
rect 9719 -202 9801 -120
rect 6154 -304 6208 -250
rect 6470 -304 6524 -250
rect 6786 -304 6840 -250
rect 7102 -304 7156 -250
rect 7418 -304 7472 -250
rect 7734 -304 7788 -250
rect 8050 -304 8104 -250
rect 8366 -304 8420 -250
rect 8682 -304 8736 -250
rect 8998 -304 9052 -250
rect 9847 -318 9929 -236
rect 5988 -1976 6042 -1922
rect 6304 -1976 6358 -1922
rect 6620 -1976 6674 -1922
rect 6936 -1976 6990 -1922
rect 7252 -1976 7306 -1922
rect 7568 -1976 7622 -1922
rect 7884 -1976 7938 -1922
rect 8200 -1976 8254 -1922
rect 8516 -1976 8570 -1922
rect 8832 -1976 8886 -1922
rect 9148 -1976 9202 -1922
rect 9847 -1990 9937 -1900
rect 6144 -2090 6198 -2036
rect 6460 -2090 6514 -2036
rect 6776 -2090 6830 -2036
rect 7092 -2090 7146 -2036
rect 7408 -2090 7462 -2036
rect 7724 -2090 7778 -2036
rect 8040 -2090 8094 -2036
rect 8356 -2090 8410 -2036
rect 8672 -2090 8726 -2036
rect 8988 -2090 9042 -2036
rect 9607 -2253 9689 -2171
<< metal2 >>
rect 9719 -120 9801 -114
rect 5988 -134 9719 -120
rect 5988 -188 5998 -134
rect 6052 -188 6314 -134
rect 6368 -188 6630 -134
rect 6684 -188 6946 -134
rect 7000 -188 7262 -134
rect 7316 -188 7578 -134
rect 7632 -188 7894 -134
rect 7948 -188 8210 -134
rect 8264 -188 8526 -134
rect 8580 -188 8842 -134
rect 8896 -188 9158 -134
rect 9212 -188 9719 -134
rect 5988 -202 9719 -188
rect 9719 -208 9801 -202
rect 9847 -236 9929 -230
rect 6144 -250 9847 -236
rect 6144 -304 6154 -250
rect 6208 -304 6470 -250
rect 6524 -304 6786 -250
rect 6840 -304 7102 -250
rect 7156 -304 7418 -250
rect 7472 -304 7734 -250
rect 7788 -304 8050 -250
rect 8104 -304 8366 -250
rect 8420 -304 8682 -250
rect 8736 -304 8998 -250
rect 9052 -304 9847 -250
rect 6144 -318 9847 -304
rect 9847 -324 9929 -318
rect 9847 -1900 9937 -1894
rect 5978 -1922 9847 -1900
rect 5978 -1976 5988 -1922
rect 6042 -1976 6304 -1922
rect 6358 -1976 6620 -1922
rect 6674 -1976 6936 -1922
rect 6990 -1976 7252 -1922
rect 7306 -1976 7568 -1922
rect 7622 -1976 7884 -1922
rect 7938 -1976 8200 -1922
rect 8254 -1976 8516 -1922
rect 8570 -1976 8832 -1922
rect 8886 -1976 9148 -1922
rect 9202 -1976 9847 -1922
rect 5978 -1990 9847 -1976
rect 9847 -1996 9937 -1990
rect 6134 -2036 9689 -2022
rect 6134 -2090 6144 -2036
rect 6198 -2090 6460 -2036
rect 6514 -2090 6776 -2036
rect 6830 -2090 7092 -2036
rect 7146 -2090 7408 -2036
rect 7462 -2090 7724 -2036
rect 7778 -2090 8040 -2036
rect 8094 -2090 8356 -2036
rect 8410 -2090 8672 -2036
rect 8726 -2090 8988 -2036
rect 9042 -2090 9689 -2036
rect 6134 -2104 9689 -2090
rect 9607 -2171 9689 -2104
rect 9607 -2259 9689 -2253
use sky130_fd_pr__pfet_g5v0d10v5_CRUJC2  XM1
timestamp 1757256347
transform 1 0 3920 0 1 -230
box -308 -362 308 362
use sky130_fd_pr__nfet_g5v0d10v5_RGPY9J  XM2
timestamp 1757256469
transform 1 0 7595 0 1 -1975
box -1781 -327 1781 327
use sky130_fd_pr__pfet_g5v0d10v5_2ZQPNU  XM3
timestamp 1757256469
transform 1 0 7605 0 1 -256
box -1809 -362 1809 362
use sky130_fd_pr__nfet_g5v0d10v5_AWMRGD  XM5
timestamp 1757256347
transform 1 0 3891 0 1 -1996
box -280 -327 280 327
<< labels >>
flabel metal1 3626 830 3826 1030 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 3636 -3030 3836 -2830 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 2992 -1188 3192 -988 0 FreeSans 256 0 0 0 input
port 3 nsew
flabel metal1 9784 -1182 9984 -982 0 FreeSans 256 0 0 0 output
port 2 nsew
<< end >>
