magic
tech sky130A
magscale 1 2
timestamp 1757299738
<< metal1 >>
rect 15126 6492 15526 6498
rect 15526 6092 26456 6492
rect 15126 6086 15526 6092
rect 18152 4354 18332 4360
rect 18332 4174 19690 4354
rect 18152 4168 18332 4174
rect 26310 4170 27414 4350
rect 14254 2588 14654 2594
rect 14654 2188 26436 2588
rect 27234 2508 27414 4170
rect 27228 2328 27234 2508
rect 27414 2328 27420 2508
rect 14254 2182 14654 2188
<< via1 >>
rect 15126 6092 15526 6492
rect 18152 4174 18332 4354
rect 14254 2188 14654 2588
rect 27234 2328 27414 2508
<< metal2 >>
rect 12875 6492 13265 6496
rect 12870 6487 15126 6492
rect 12870 6097 12875 6487
rect 13265 6097 15126 6487
rect 12870 6092 15126 6097
rect 15526 6092 15532 6492
rect 12875 6088 13265 6092
rect 18146 4174 18152 4354
rect 18332 4174 18338 4354
rect 11257 2588 11647 2592
rect 11252 2583 14254 2588
rect 11252 2193 11257 2583
rect 11647 2193 14254 2583
rect 11252 2188 14254 2193
rect 14654 2188 14660 2588
rect 11257 2184 11647 2188
rect 18152 1581 18332 4174
rect 27234 2508 27414 2514
rect 27234 1977 27414 2328
rect 27230 1807 27239 1977
rect 27409 1807 27418 1977
rect 27234 1802 27414 1807
rect 18152 1411 18157 1581
rect 18327 1411 18332 1581
rect 18152 1406 18332 1411
rect 18157 1402 18327 1406
<< via2 >>
rect 12875 6097 13265 6487
rect 11257 2193 11647 2583
rect 27239 1807 27409 1977
rect 18157 1411 18327 1581
<< metal3 >>
rect 4577 6492 4975 6497
rect 4576 6491 13270 6492
rect 4576 6093 4577 6491
rect 4975 6487 13270 6491
rect 4975 6097 12875 6487
rect 13265 6097 13270 6487
rect 4975 6093 13270 6097
rect 4576 6092 13270 6093
rect 4577 6087 4975 6092
rect 9789 2588 10187 2593
rect 9788 2587 11652 2588
rect 9788 2189 9789 2587
rect 10187 2583 11652 2587
rect 10187 2193 11257 2583
rect 11647 2193 11652 2583
rect 10187 2189 11652 2193
rect 9788 2188 11652 2189
rect 9789 2183 10187 2188
rect 27234 1977 27414 1982
rect 27234 1807 27239 1977
rect 27409 1807 27414 1977
rect 23371 1586 23549 1591
rect 18152 1585 23550 1586
rect 18152 1581 23371 1585
rect 18152 1411 18157 1581
rect 18327 1411 23371 1581
rect 18152 1407 23371 1411
rect 23549 1407 23550 1585
rect 27234 1531 27414 1807
rect 18152 1406 23550 1407
rect 23371 1401 23549 1406
rect 27229 1353 27235 1531
rect 27413 1353 27419 1531
rect 27234 1352 27414 1353
<< via3 >>
rect 4577 6093 4975 6491
rect 9789 2189 10187 2587
rect 23371 1407 23549 1585
rect 27235 1353 27413 1531
<< metal4 >>
rect 3006 44776 3066 45152
rect 3558 44776 3618 45152
rect 4110 44776 4170 45152
rect 4662 44776 4722 45152
rect 5214 44776 5274 45152
rect 5766 44776 5826 45152
rect 6318 44776 6378 45152
rect 6870 44776 6930 45152
rect 7422 44776 7482 45152
rect 7974 44776 8034 45152
rect 8526 44776 8586 45152
rect 9078 44776 9138 45152
rect 9630 45062 9690 45152
rect 9622 44952 9690 45062
rect 9622 44776 9682 44952
rect 10182 44776 10242 45152
rect 10734 44776 10794 45152
rect 11286 44776 11346 45152
rect 11838 44776 11898 45152
rect 12390 44776 12450 45152
rect 12942 44776 13002 45152
rect 13494 44776 13554 45152
rect 14046 44776 14106 45152
rect 14598 44776 14658 45152
rect 15150 44776 15210 45152
rect 15702 44776 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 3004 44396 15800 44776
rect 3592 6492 3992 44138
rect 3592 6491 4976 6492
rect 3592 6093 4577 6491
rect 4975 6093 4976 6491
rect 3592 6092 4976 6093
rect 3592 986 3992 6092
rect 6000 2588 6400 44396
rect 6000 2587 10188 2588
rect 6000 2189 9789 2587
rect 10187 2189 10188 2587
rect 6000 2188 10188 2189
rect 6000 990 6400 2188
rect 23370 1585 23550 1586
rect 23370 1407 23371 1585
rect 23549 1407 23550 1585
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 1407
rect 27234 1531 27414 1532
rect 27234 1353 27235 1531
rect 27413 1353 27414 1531
rect 27234 0 27414 1353
use double_inverter  double_inverter_0
timestamp 1757295524
transform 1 0 16510 0 1 5342
box 2992 -3030 9984 1030
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 6000 990 6400 44142 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 3592 986 3992 44138 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
